library ieee;
use ieee.std_logic_1164.all;

entity logic_unit is
    port(
        a  : in  std_logic_vector(31 downto 0);
        b  : in  std_logic_vector(31 downto 0);
        op : in  std_logic_vector(1 downto 0);
        r  : out std_logic_vector(31 downto 0)
    );
end logic_unit;

architecture synth of logic_unit is
BEGIN
  
  r <= (a NOR b) WHEN op = "00" ELSE
	(a AND b) WHEN op = "01" ELSE
	(a OR b) WHEN op = "10" ELSE
	(a XNOR b) WHEN op = "11" ELSE
	(others => '0');

end synth;
